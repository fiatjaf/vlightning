module vlightning
